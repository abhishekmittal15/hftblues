package TestBench;

// Imports 
import LFSR::*;




endpackage: TestBench
