package C_imports;

	import "BDPI" function ActionValue #(Bit #(32)) get_packet();

endpackage: C_imports
