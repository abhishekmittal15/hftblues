/* package declaration */ 

