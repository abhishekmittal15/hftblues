package deepthought;

module DeepThought;

    rule RuleName(Cond);
        
    endrule

endmodule
