package c_imports;

import "BDPI" function ActionValue #(Int#(32)) open_file();

import "BDPI" function ActionValue #(Int#(32)) read_ints();

import "BDPI" function ActionValue #(Int#(32)) close_file();

endpackage: c_imports